`include "parallel_prefix.v"

module cla_adder(a, b, sum, c);

    input [31:0] a, b;
    output [31:0] sum;
    output c;
    
    wire [63:0] kpg, kpg1, kpg2, kpg3, kpg4, kpg5;
    wire [31:0] carry;

    assign kpg[0] = a[0];
    assign kpg[1] = b[0];
    assign kpg[2] = a[1];
    assign kpg[3] = b[1];
    assign kpg[4] = a[2];
    assign kpg[5] = b[2];
    assign kpg[6] = a[3];
    assign kpg[7] = b[3];
    assign kpg[8] = a[4];
    assign kpg[9] = b[4];
    assign kpg[10] = a[5];
    assign kpg[11] = b[5];
    assign kpg[12] = a[6];
    assign kpg[13] = b[6];
    assign kpg[14] = a[7];
    assign kpg[15] = b[7];
    assign kpg[16] = a[8];
    assign kpg[17] = b[8];
    assign kpg[18] = a[9];
    assign kpg[19] = b[9];
    assign kpg[20] = a[10];
    assign kpg[21] = b[10];
    assign kpg[22] = a[11];
    assign kpg[23] = b[11];
    assign kpg[24] = a[12];
    assign kpg[25] = b[12];
    assign kpg[26] = a[13];
    assign kpg[27] = b[13];
    assign kpg[28] = a[14];
    assign kpg[29] = b[14];
    assign kpg[30] = a[15];
    assign kpg[31] = b[15];
    assign kpg[32] = a[16];
    assign kpg[33] = b[16];
    assign kpg[34] = a[17];
    assign kpg[35] = b[17];
    assign kpg[36] = a[18];
    assign kpg[37] = b[18];
    assign kpg[38] = a[19];
    assign kpg[39] = b[19];
    assign kpg[40] = a[20];
    assign kpg[41] = b[20];
    assign kpg[42] = a[21];
    assign kpg[43] = b[21];
    assign kpg[44] = a[22];
    assign kpg[45] = b[22];
    assign kpg[46] = a[23];
    assign kpg[47] = b[23];
    assign kpg[48] = a[24];
    assign kpg[49] = b[24];
    assign kpg[50] = a[25];
    assign kpg[51] = b[25];
    assign kpg[52] = a[26];
    assign kpg[53] = b[26];
    assign kpg[54] = a[27];
    assign kpg[55] = b[27];
    assign kpg[56] = a[28];
    assign kpg[57] = b[28];
    assign kpg[58] = a[29];
    assign kpg[59] = b[29];
    assign kpg[60] = a[30];
    assign kpg[61] = b[30];
    assign kpg[62] = a[31];
    assign kpg[63] = b[31];


    parallelprefix p0(kpg[1:0], 2'b00, kpg1[1:0]);
    parallelprefix p1(kpg[3:2], kpg1[1:0], kpg1[3:2]);
    parallelprefix p2(kpg[5:4], kpg1[3:2], kpg1[5:4]);
    parallelprefix p3(kpg[7:6], kpg1[5:4], kpg1[7:6]);
    parallelprefix p4(kpg[9:8], kpg1[7:6], kpg1[9:8]);
    parallelprefix p5(kpg[11:10], kpg1[9:8], kpg1[11:10]);
    parallelprefix p6(kpg[13:12], kpg1[11:10], kpg1[13:12]);
    parallelprefix p7(kpg[15:14], kpg1[13:12], kpg1[15:14]);
    parallelprefix p8(kpg[17:16], kpg1[15:14], kpg1[17:16]);
    parallelprefix p9(kpg[19:18], kpg1[17:16], kpg1[19:18]);
    parallelprefix p10(kpg[21:20], kpg1[19:18], kpg1[21:20]);
    parallelprefix p11(kpg[23:22], kpg1[21:20], kpg1[23:22]);
    parallelprefix p12(kpg[25:24], kpg1[23:22], kpg1[25:24]);
    parallelprefix p13(kpg[27:26], kpg1[25:24], kpg1[27:26]);
    parallelprefix p14(kpg[29:28], kpg1[27:26], kpg1[29:28]);
    parallelprefix p15(kpg[31:30], kpg1[29:28], kpg1[31:30]);
    parallelprefix p16(kpg[33:32], kpg1[31:30], kpg1[33:32]);
    parallelprefix p17(kpg[35:34], kpg1[33:32], kpg1[35:34]);
    parallelprefix p18(kpg[37:36], kpg1[35:34], kpg1[37:36]);
    parallelprefix p19(kpg[39:38], kpg1[37:36], kpg1[39:38]);
    parallelprefix p20(kpg[41:40], kpg1[39:38], kpg1[41:40]);
    parallelprefix p21(kpg[43:42], kpg1[41:40], kpg1[43:42]);
    parallelprefix p22(kpg[45:44], kpg1[43:42], kpg1[45:44]);
    parallelprefix p23(kpg[47:46], kpg1[45:44], kpg1[47:46]);
    parallelprefix p24(kpg[49:48], kpg1[47:46], kpg1[49:48]);
    parallelprefix p25(kpg[51:50], kpg1[49:48], kpg1[51:50]);
    parallelprefix p26(kpg[53:52], kpg1[51:50], kpg1[53:52]);
    parallelprefix p27(kpg[55:54], kpg1[53:52], kpg1[55:54]);
    parallelprefix p28(kpg[57:56], kpg1[55:54], kpg1[57:56]);
    parallelprefix p29(kpg[59:58], kpg1[57:56], kpg1[59:58]);
    parallelprefix p30(kpg[61:60], kpg1[59:58], kpg1[61:60]);
    parallelprefix p31(kpg[63:62], kpg1[61:60], kpg1[63:62]);


    parallelprefix p32(kpg1[1:0], 2'b00, kpg2[1:0]);
    parallelprefix p33(kpg1[3:2], 2'b00, kpg2[3:2]);
    parallelprefix p34(kpg1[5:4], kpg2[3:2], kpg2[5:4]);
    parallelprefix p35(kpg1[7:6], kpg2[5:4], kpg2[7:6]);
    parallelprefix p36(kpg1[9:8], kpg2[7:6], kpg2[9:8]);
    parallelprefix p37(kpg1[11:10], kpg2[9:8], kpg2[11:10]);
    parallelprefix p38(kpg1[13:12], kpg2[11:10], kpg2[13:12]);
    parallelprefix p39(kpg1[15:14], kpg2[13:12], kpg2[15:14]);
    parallelprefix p40(kpg1[17:16], kpg2[15:14], kpg2[17:16]);
    parallelprefix p41(kpg1[19:18], kpg2[17:16], kpg2[19:18]);
    parallelprefix p42(kpg1[21:20], kpg2[19:18], kpg2[21:20]);
    parallelprefix p43(kpg1[23:22], kpg2[21:20], kpg2[23:22]);
    parallelprefix p44(kpg1[25:24], kpg2[23:22], kpg2[25:24]);
    parallelprefix p45(kpg1[27:26], kpg2[25:24], kpg2[27:26]);
    parallelprefix p46(kpg1[29:28], kpg2[27:26], kpg2[29:28]);
    parallelprefix p47(kpg1[31:30], kpg2[29:28], kpg2[31:30]);
    parallelprefix p48(kpg1[33:32], kpg2[31:30], kpg2[33:32]);
    parallelprefix p49(kpg1[35:34], kpg2[33:32], kpg2[35:34]);
    parallelprefix p50(kpg1[37:36], kpg2[35:34], kpg2[37:36]);
    parallelprefix p51(kpg1[39:38], kpg2[37:36], kpg2[39:38]);
    parallelprefix p52(kpg1[41:40], kpg2[39:38], kpg2[41:40]);
    parallelprefix p53(kpg1[43:42], kpg2[41:40], kpg2[43:42]);
    parallelprefix p54(kpg1[45:44], kpg2[43:42], kpg2[45:44]);
    parallelprefix p55(kpg1[47:46], kpg2[45:44], kpg2[47:46]);
    parallelprefix p56(kpg1[49:48], kpg2[47:46], kpg2[49:48]);
    parallelprefix p57(kpg1[51:50], kpg2[49:48], kpg2[51:50]);
    parallelprefix p58(kpg1[53:52], kpg2[51:50], kpg2[53:52]);
    parallelprefix p59(kpg1[55:54], kpg2[53:52], kpg2[55:54]);
    parallelprefix p60(kpg1[57:56], kpg2[55:54], kpg2[57:56]);
    parallelprefix p61(kpg1[59:58], kpg2[57:56], kpg2[59:58]);
    parallelprefix p62(kpg1[61:60], kpg2[59:58], kpg2[61:60]);
    parallelprefix p63(kpg1[63:62], kpg2[61:60], kpg2[63:62]);



    parallelprefix p64(kpg2[1:0], 2'b00, kpg3[1:0]);
    parallelprefix p65(kpg2[3:2], 2'b00, kpg3[3:2]);
    parallelprefix p66(kpg2[5:4], 2'b00, kpg3[5:4]);
    parallelprefix p67(kpg2[7:6], 2'b00, kpg3[7:6]);
    parallelprefix p68(kpg2[9:8], kpg3[7:6], kpg3[9:8]);
    parallelprefix p69(kpg2[11:10], kpg3[9:8], kpg3[11:10]);
    parallelprefix p70(kpg2[13:12], kpg3[11:10], kpg3[13:12]);
    parallelprefix p71(kpg2[15:14], kpg3[13:12], kpg3[15:14]);
    parallelprefix p72(kpg2[17:16], kpg3[15:14], kpg3[17:16]);
    parallelprefix p73(kpg2[19:18], kpg3[17:16], kpg3[19:18]);
    parallelprefix p74(kpg2[21:20], kpg3[19:18], kpg3[21:20]);
    parallelprefix p75(kpg2[23:22], kpg3[21:20], kpg3[23:22]);
    parallelprefix p76(kpg2[25:24], kpg3[23:22], kpg3[25:24]);
    parallelprefix p77(kpg2[27:26], kpg3[25:24], kpg3[27:26]);
    parallelprefix p78(kpg2[29:28], kpg3[27:26], kpg3[29:28]);
    parallelprefix p79(kpg2[31:30], kpg3[29:28], kpg3[31:30]);
    parallelprefix p80(kpg2[33:32], kpg3[31:30], kpg3[33:32]);
    parallelprefix p81(kpg2[35:34], kpg3[33:32], kpg3[35:34]);
    parallelprefix p82(kpg2[37:36], kpg3[35:34], kpg3[37:36]);
    parallelprefix p83(kpg2[39:38], kpg3[37:36], kpg3[39:38]);
    parallelprefix p84(kpg2[41:40], kpg3[39:38], kpg3[41:40]);
    parallelprefix p85(kpg2[43:42], kpg3[41:40], kpg3[43:42]);
    parallelprefix p86(kpg2[45:44], kpg3[43:42], kpg3[45:44]);
    parallelprefix p87(kpg2[47:46], kpg3[45:44], kpg3[47:46]);
    parallelprefix p88(kpg2[49:48], kpg3[47:46], kpg3[49:48]);
    parallelprefix p89(kpg2[51:50], kpg3[49:48], kpg3[51:50]);
    parallelprefix p90(kpg2[53:52], kpg3[51:50], kpg3[53:52]);
    parallelprefix p91(kpg2[55:54], kpg3[53:52], kpg3[55:54]);
    parallelprefix p92(kpg2[57:56], kpg3[55:54], kpg3[57:56]);
    parallelprefix p93(kpg2[59:58], kpg3[57:56], kpg3[59:58]);
    parallelprefix p94(kpg2[61:60], kpg3[59:58], kpg3[61:60]);
    parallelprefix p95(kpg2[63:62], kpg3[61:60], kpg3[63:62]);


    parallelprefix p96(kpg3[3:2], 2'b00, kpg4[3:2]);
    parallelprefix p97(kpg3[3:2], 2'b00, kpg4[3:2]);
    parallelprefix p98(kpg3[5:4], 2'b00, kpg4[5:4]);
    parallelprefix p99(kpg3[7:6], 2'b00, kpg4[7:6]);
    parallelprefix p100(kpg3[9:8], 2'b00, kpg4[9:8]);
    parallelprefix p101(kpg3[11:10], 2'b00, kpg4[11:10]);
    parallelprefix p102(kpg3[13:12], 2'b00, kpg4[13:12]);
    parallelprefix p103(kpg3[15:14], 2'b00, kpg4[15:14]);
    parallelprefix p104(kpg3[17:16], kpg4[15:14], kpg4[17:16]);
    parallelprefix p105(kpg3[19:18], kpg4[17:16], kpg4[19:18]);
    parallelprefix p106(kpg3[21:20], kpg4[19:18], kpg4[21:20]);
    parallelprefix p107(kpg3[23:22], kpg4[21:20], kpg4[23:22]);
    parallelprefix p108(kpg3[25:24], kpg4[23:22], kpg4[25:24]);
    parallelprefix p109(kpg3[27:26], kpg4[25:24], kpg4[27:26]);
    parallelprefix p110(kpg3[29:28], kpg4[27:26], kpg4[29:28]);
    parallelprefix p111(kpg3[31:30], kpg4[29:28], kpg4[31:30]);
    parallelprefix p112(kpg3[33:32], kpg4[31:30], kpg4[33:32]);
    parallelprefix p113(kpg3[35:34], kpg4[33:32], kpg4[35:34]);
    parallelprefix p114(kpg3[37:36], kpg4[35:34], kpg4[37:36]);
    parallelprefix p115(kpg3[39:38], kpg4[37:36], kpg4[39:38]);
    parallelprefix p116(kpg3[41:40], kpg4[39:38], kpg4[41:40]);
    parallelprefix p117(kpg3[43:42], kpg4[41:40], kpg4[43:42]);
    parallelprefix p118(kpg3[45:44], kpg4[43:42], kpg4[45:44]);
    parallelprefix p119(kpg3[47:46], kpg4[45:44], kpg4[47:46]);
    parallelprefix p120(kpg3[49:48], kpg4[47:46], kpg4[49:48]);
    parallelprefix p121(kpg3[51:50], kpg4[49:48], kpg4[51:50]);
    parallelprefix p122(kpg3[53:52], kpg4[51:50], kpg4[53:52]);
    parallelprefix p123(kpg3[55:54], kpg4[53:52], kpg4[55:54]);
    parallelprefix p124(kpg3[57:56], kpg4[55:54], kpg4[57:56]);
    parallelprefix p125(kpg3[59:58], kpg4[57:56], kpg4[59:58]);
    parallelprefix p126(kpg3[61:60], kpg4[59:58], kpg4[61:60]);
    parallelprefix p127(kpg3[63:62], kpg4[61:60], kpg4[63:62]);

    parallelprefix p128(kpg4[1:0], 2'b00, kpg5[1:0]);
    parallelprefix p129(kpg4[3:2], 2'b00, kpg5[3:2]);
    parallelprefix p130(kpg4[5:4], 2'b00, kpg5[5:4]);
    parallelprefix p131(kpg4[7:6], 2'b00, kpg5[7:6]);
    parallelprefix p132(kpg4[9:8], 2'b00, kpg5[9:8]);
    parallelprefix p133(kpg4[11:10], 2'b00, kpg5[11:10]);
    parallelprefix p134(kpg4[13:12], 2'b00, kpg5[13:12]);
    parallelprefix p135(kpg4[15:14], 2'b00, kpg5[15:14]);
    parallelprefix p136(kpg4[17:16], 2'b00, kpg5[17:16]);
    parallelprefix p137(kpg4[19:18], 2'b00, kpg5[19:18]);
    parallelprefix p138(kpg4[21:20], 2'b00, kpg5[21:20]);
    parallelprefix p139(kpg4[23:22], 2'b00, kpg5[23:22]);
    parallelprefix p140(kpg4[25:24], 2'b00, kpg5[25:24]);
    parallelprefix p141(kpg4[27:26], 2'b00, kpg5[27:26]);
    parallelprefix p142(kpg4[29:28], 2'b00, kpg5[29:28]);
    parallelprefix p143(kpg4[31:30], 2'b00, kpg5[31:30]);
    parallelprefix p144(kpg4[33:32], kpg5[31:30], kpg5[33:32]);
    parallelprefix p145(kpg4[35:34], kpg5[33:32], kpg5[35:34]);
    parallelprefix p146(kpg4[37:36], kpg5[35:34], kpg5[37:36]);
    parallelprefix p147(kpg4[39:38], kpg5[37:36], kpg5[39:38]);
    parallelprefix p148(kpg4[41:40], kpg5[39:38], kpg5[41:40]);
    parallelprefix p149(kpg4[43:42], kpg5[41:40], kpg5[43:42]);
    parallelprefix p150(kpg4[45:44], kpg5[43:42], kpg5[45:44]);
    parallelprefix p151(kpg4[47:46], kpg5[45:44], kpg5[47:46]);
    parallelprefix p152(kpg4[49:48], kpg5[47:46], kpg5[49:48]);
    parallelprefix p153(kpg4[51:50], kpg5[49:48], kpg5[51:50]);
    parallelprefix p154(kpg4[53:52], kpg5[51:50], kpg5[53:52]);
    parallelprefix p155(kpg4[55:54], kpg5[53:52], kpg5[55:54]);
    parallelprefix p156(kpg4[57:56], kpg5[55:54], kpg5[57:56]);
    parallelprefix p157(kpg4[59:58], kpg5[57:56], kpg5[59:58]);
    parallelprefix p158(kpg4[61:60], kpg5[59:58], kpg5[61:60]);
    parallelprefix p159(kpg4[63:62], kpg5[61:60], kpg5[63:62]);


    assign carry[0] = kpg5[1];
    assign carry[1] = kpg5[3];
    assign carry[2] = kpg5[5];
    assign carry[3] = kpg5[7];
    assign carry[4] = kpg5[9];
    assign carry[5] = kpg5[11];
    assign carry[6] = kpg5[13];
    assign carry[7] = kpg5[15];
    assign carry[8] = kpg5[17];
    assign carry[9] = kpg5[19];
    assign carry[10] = kpg5[21];
    assign carry[11] = kpg5[23];
    assign carry[12] = kpg5[25];
    assign carry[13] = kpg5[27];
    assign carry[14] = kpg5[29];
    assign carry[15] = kpg5[31];
    assign carry[16] = kpg5[33];
    assign carry[17] = kpg5[35];
    assign carry[18] = kpg5[37];
    assign carry[19] = kpg5[39];
    assign carry[20] = kpg5[41];
    assign carry[21] = kpg5[43];
    assign carry[22] = kpg5[45];
    assign carry[23] = kpg5[47];
    assign carry[24] = kpg5[49];
    assign carry[25] = kpg5[51];
    assign carry[26] = kpg5[53];
    assign carry[27] = kpg5[55];
    assign carry[28] = kpg5[57];
    assign carry[29] = kpg5[59];
    assign carry[30] = kpg5[61];
    assign carry[31] = kpg5[63];

    assign sum[0] = a[0] ^ b[0];
    assign sum[1] = a[1] ^ b[1] ^ carry[0];
    assign sum[2] = a[2] ^ b[2] ^ carry[1];
    assign sum[3] = a[3] ^ b[3] ^ carry[2];
    assign sum[4] = a[4] ^ b[4] ^ carry[3];
    assign sum[5] = a[5] ^ b[5] ^ carry[4];
    assign sum[6] = a[6] ^ b[6] ^ carry[5];
    assign sum[7] = a[7] ^ b[7] ^ carry[6];
    assign sum[8] = a[8] ^ b[8] ^ carry[7];
    assign sum[9] = a[9] ^ b[9] ^ carry[8];
    assign sum[10] = a[10] ^ b[10] ^ carry[9];
    assign sum[11] = a[11] ^ b[11] ^ carry[10];
    assign sum[12] = a[12] ^ b[12] ^ carry[11];
    assign sum[13] = a[13] ^ b[13] ^ carry[12];
    assign sum[14] = a[14] ^ b[14] ^ carry[13];
    assign sum[15] = a[15] ^ b[15] ^ carry[14];
    assign sum[16] = a[16] ^ b[16] ^ carry[15];
    assign sum[17] = a[17] ^ b[17] ^ carry[16];
    assign sum[18] = a[18] ^ b[18] ^ carry[17];
    assign sum[19] = a[19] ^ b[19] ^ carry[18];
    assign sum[20] = a[20] ^ b[20] ^ carry[19];
    assign sum[21] = a[21] ^ b[21] ^ carry[20];
    assign sum[22] = a[22] ^ b[22] ^ carry[21];
    assign sum[23] = a[23] ^ b[23] ^ carry[22];
    assign sum[24] = a[24] ^ b[24] ^ carry[23];
    assign sum[25] = a[25] ^ b[25] ^ carry[24];
    assign sum[26] = a[26] ^ b[26] ^ carry[25];
    assign sum[27] = a[27] ^ b[27] ^ carry[26];
    assign sum[28] = a[28] ^ b[28] ^ carry[27];
    assign sum[29] = a[29] ^ b[29] ^ carry[28];
    assign sum[30] = a[30] ^ b[30] ^ carry[29];
    assign sum[31] = a[31] ^ b[31] ^ carry[30];
    assign c = carry[31];

endmodule
