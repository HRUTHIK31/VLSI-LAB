magic
tech scmos
timestamp 1597289998
<< nwell >>
rect -52 7 -10 18
rect -1 7 45 18
<< polysilicon >>
rect -42 16 -39 20
rect -25 16 -22 20
rect 21 16 24 20
rect -42 -17 -39 9
rect -25 -17 -22 9
rect 21 -2 24 9
rect -7 -8 24 -2
rect 21 -17 24 -8
rect -42 -26 -39 -24
rect -25 -26 -22 -24
rect 21 -26 24 -24
<< ndiffusion >>
rect -44 -24 -42 -17
rect -39 -24 -25 -17
rect -22 -24 -19 -17
rect 8 -24 21 -17
rect 24 -24 36 -17
<< pdiffusion >>
rect -44 9 -42 16
rect -39 9 -36 16
rect -28 9 -25 16
rect -22 9 -18 16
rect 9 9 21 16
rect 24 9 36 16
<< metal1 >>
rect -52 22 -42 29
rect -35 22 -25 29
rect -18 22 -5 29
rect 2 22 15 29
rect 22 22 32 29
rect 39 22 45 29
rect -50 16 -44 22
rect -18 16 -12 22
rect 1 16 9 22
rect -36 1 -28 9
rect -36 -7 -13 1
rect -19 -17 -13 -7
rect 36 -17 43 9
rect -50 -28 -44 -24
rect 1 -28 8 -24
rect -50 -36 -41 -28
rect -34 -36 -23 -28
rect -16 -36 -7 -28
rect 0 -36 17 -28
rect 24 -36 36 -28
rect 43 -36 49 -28
<< ntransistor >>
rect -42 -24 -39 -17
rect -25 -24 -22 -17
rect 21 -24 24 -17
<< ptransistor >>
rect -42 9 -39 16
rect -25 9 -22 16
rect 21 9 24 16
<< polycontact >>
rect -13 -8 -7 -2
<< ndcontact >>
rect -50 -24 -44 -17
rect -19 -24 -13 -17
rect 1 -24 8 -17
rect 36 -24 43 -17
<< pdcontact >>
rect -50 9 -44 16
rect -36 9 -28 16
rect -18 9 -12 16
rect 1 9 9 16
rect 36 9 43 16
<< psubstratepcontact >>
rect -41 -36 -34 -28
rect -23 -36 -16 -28
rect -7 -36 0 -28
rect 17 -36 24 -28
rect 36 -36 43 -28
<< nsubstratencontact >>
rect -42 22 -35 29
rect -25 22 -18 29
rect -5 22 2 29
rect 15 22 22 29
rect 32 22 39 29
<< labels >>
rlabel metal1 -48 24 -48 24 4 vdd
rlabel metal1 -47 -33 -47 -33 2 gnd
rlabel polysilicon -41 -12 -41 -12 1 a
rlabel polysilicon -24 -12 -24 -12 1 b
rlabel metal1 39 -11 39 -11 1 y
<< end >>
